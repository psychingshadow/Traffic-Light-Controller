module Traffic_Light_Controller_TB;
    reg clk, reset;
    wire [2 : 0] light_M1;
    wire [2 : 0] light_S;
    wire [2 : 0] light_MT;
    wire [2 : 0] light_M2;

Traffic_Light_Controller TLC(.clk(clk), .reset(reset), .light_M1(light_M1), .light_S(light_S), .light_M2(light_M2), .light_MT(light_MT));

    initial
	begin
    	    clk = 1'b0;
    	    forever #(1000000000/2) clk = ~clk;
	end

    initial
	begin
            reset = 0;
            #1000000000;
            reset = 1;
            #1000000000;
            reset = 0;
   	end
endmodule